library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top_module is
end top_module;

architecture Behavioral of top_module is

begin


end Behavioral;

